module InstructionMemory
(
    output  logic [31:0] instruction_data_o,
    input   logic [31:0] instruction_address_i
);

    logic [31:0] instruction [63:0];

    initial 
    begin
        $readmesh("L_S_type.txt", instruction);
    end

    always_comb
    begin
        instruction_data_o = instruction[instruction_address_i[31:2]];
    end

endmodule